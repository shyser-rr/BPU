module extend_unit (
    input logic [2:0] imm_src
);

endmodule